module seg (
    ports
);
    
endmodule